typedef enum logic[3:0] {
    DECODE,
    ALIGN,
    OPERATE,
    NORMALIZE,
    WRITEBACK
} state_t;

typedef enum logic[3:0] { 
    OVERFLOW,
    UNDERFLOW,
    EXACT,
    INEXACT
} status_t;

module FPU(
    input  logic        clock_100Khz,
    input  logic        reset,      // assíncrono ativo-baixo
    input  logic [31:0] Op_A_in,
    input  logic [31:0] Op_B_in,
    output logic [31:0] data_out,
    output status_t     status_out
);

    state_t EA, PE;

    // sinais auxiliares
    logic sign_A, sign_B, carry, compare;
    logic done_decode, done_align, done_operate, done_normalize, done_writeback;

    // campos de mantissa e expoente
    logic [21:0] mant_A, mant_B, mant_SHIFT, mant_TMP, mant_A_tmp, mant_B_tmp;
    logic [9:0]  exp_A, exp_B, exp_TMP, exp_A_tmp, exp_B_tmp;
    logic [9:0]  diff_Exponent;

    // FSM sequencial
    always_ff @(posedge clock_100Khz or negedge reset) begin
        if (!reset) begin
            EA             <= DECODE;
            // reset flags e regs
            done_decode    <= 0; done_align <= 0; done_operate <= 0;
            done_normalize <= 0; done_writeback <= 0;
            mant_A         <= 0; mant_B <= 0; mant_SHIFT <= 0; mant_TMP<=0;
            exp_A          <= 0; exp_B<=0; exp_TMP<=0;
            sign_A         <= 0; sign_B<=0;
            data_out       <= 0; status_out <= EXACT;
            diff_Exponent  <= 0;
        end else begin
            EA <= PE;
            // ações de cada estado
            case (EA)
                DECODE: begin
                    // Prepara A e B e difere expoente
                    mant_A      <= mant_A_tmp;
                    exp_A       <= exp_A_tmp;
                    sign_A      <= compare ? Op_A_in[31] : Op_B_in[31];
                    mant_B      <= mant_B_tmp;
                    exp_B       <= exp_B_tmp;
                    sign_B      <= compare ? Op_B_in[31] : Op_A_in[31];
                    diff_Exponent<= exp_A_tmp - exp_B_tmp;
                    done_decode <= 1;
                end

                ALIGN: begin
                    // Repete shift até diff=0
                    if (diff_Exponent > 0) begin
                        mant_B        <= mant_B >> 1;
                        diff_Exponent <= diff_Exponent - 1;
                    end else begin
                        done_align    <= 1;
                        mant_SHIFT    <= mant_B;
                    end
                end

                OPERATE: begin
                    // usa mant_SHIFT já alinhado
                    if (sign_A == sign_B) {carry, mant_TMP} <= mant_A + mant_SHIFT;
                    else                  mant_TMP         <= mant_A - mant_SHIFT;
                    exp_TMP <= exp_A;
                    if (carry) begin
                        mant_TMP <= mant_TMP >> 1;
                        exp_TMP  <= exp_TMP + 1;
                    end
                    done_operate <= 1;
                end

                NORMALIZE: begin
                    // shift left até MSB em bit21
                    if (!done_normalize) begin
                        if (!mant_TMP[21]) begin
                            mant_TMP <= mant_TMP << 1;
                            exp_TMP  <= exp_TMP - 1;
                        end else begin
                            done_normalize <= 1;
                        end
                    end
                end

                WRITEBACK: begin
                    data_out       <= {sign_A, exp_TMP, mant_TMP[20:0]};
                    if      (exp_TMP == 0)            status_out <= UNDERFLOW;
                    else if (exp_TMP == 10'd1023)     status_out <= OVERFLOW;
                    else if (mant_TMP[20:0] == 0)     status_out <= INEXACT;
                    else                               status_out <= EXACT;
                    done_writeback <= 1;
                end
            endcase
        end
    end

    // FSM combinacional
    always_comb begin
        PE = EA;
        case (EA)
            DECODE:    if (done_decode)    PE = ALIGN;
            ALIGN:     if (done_align)     PE = OPERATE;
            OPERATE:   if (done_operate)   PE = NORMALIZE;
            NORMALIZE: if (done_normalize) PE = WRITEBACK;
            WRITEBACK: if (done_writeback) PE = DECODE;
            default:   PE = DECODE;
        endcase
    end

    // separação de campos
    always_comb begin
        compare    = (Op_A_in[30:21] >= Op_B_in[30:21]);
        mant_A_tmp = compare ? {1'b1, Op_A_in[20:0]} : {1'b1, Op_B_in[20:0]};
        exp_A_tmp  = compare ? Op_A_in[30:21]       : Op_B_in[30:21];
        mant_B_tmp = compare ? {1'b1, Op_B_in[20:0]} : {1'b1, Op_A_in[20:0]};
        exp_B_tmp  = compare ? Op_B_in[30:21]       : Op_A_in[30:21];
    end

endmodule
